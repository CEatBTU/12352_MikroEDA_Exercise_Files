library IEEE;
use IEEE.std_logic_1164.all; -- import std_logic types
use IEEE.numeric_std.all; -- for type conversion to_unsigned

--library STD;
--use STD.textio.all;

--------------------------------------------------------------------------------
--!@file: mult_rtl.vhd
--!@brief: this is a simple multiplier description (generic) and iterativ
--!...
--
--!@author: Tobias Koal(TK)
--!@revision info :
-- last modification by tkoal(TK)
-- Mon Apr 13 14:27:49 CEST 2015
--------------------------------------------------------------------------------

-- entity description

entity mult_rtl is
port(
);
end entity;

-- architecture description

architecture behave of mult_rtl is


begin

end behave;

